library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity D_flip_flop is
    Port (
        DIN : in STD_LOGIC;
        CLK : in STD_LOGIC;
        Q : out STD_LOGIC
    );
end D_flip_flop;

architecture Behavioral of D_flip_flop is
    signal Q_int : STD_LOGIC;
begin
    process (CLK)
    begin
        if rising_edge(CLK) then
            Q_int <= DIN; -- Update Q on rising edge of CLK
        end if;
    end process;

    -- Output Q
    Q <= Q_int;
end Behavioral;