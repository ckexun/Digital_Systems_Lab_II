module counter10(
input clk,
input clrn,
input load,
input [3:0] D,
input en,
output Co,
output reg[3:0]Q
);

always@(posedge clk)
		begin 
		if(clrn== 1)
			begin 
			Q = 0;
			end
		else if(load == 1)
			begin 
			Q = D;
			end 
		else if(en == 0)
			begin
			Q = Q;
			end
		else if(en == 1)
			begin 
			if(Q == 9)
				Q = 0;
			else
				Q = Q + 1;
			end 
		end
		assign Co = Q[3] & Q[0] & en;
 endmodule 