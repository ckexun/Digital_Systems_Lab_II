module lab08_1 (
    input clrn, clk, Ldn, Sh, Di, D3, D2, D1, D0,
    output reg Q3, Q2, Q1, Q0
);

reg [3:0] tmp;

always @(posedge clk or posedge clrn) begin
    if (clrn) begin
        tmp <= 4'b0000; // �M���Ȧs��
    end else if (Ldn) begin
        tmp <= {D3, D2, D1, D0}; // �ñ���J���J�Ȧs��
    end
end

always @(*) begin
    case ({Ldn, Sh})
        2'b10: begin // ��XD3~D0�A�h�u����JD3~D0�����J���(���J)
            Q3 = tmp[3];
            Q2 = tmp[2];
            Q1 = tmp[1];
            Q0 = tmp[0];
        end
        2'b01: begin // ��XDi,Q3~Q1�ADi,Q3~Q1���e�ſ�X(����)
            Q3 = Di;
            Q2 = tmp[2];
            Q1 = tmp[1];
            Q0 = tmp[0];
        end
        default: begin // ��XQ3~Q0�AQ3~Q0����X�^��(����)
            Q3 = tmp[3];
            Q2 = tmp[2];
            Q1 = tmp[1];
            Q0 = tmp[0];
        end
    endcase
end

endmodule
