library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity lab13_G09 is
    Port ( clk   : in  STD_LOGIC;
           hex0  : out STD_LOGIC_VECTOR (7 downto 0);
           hex1  : out STD_LOGIC_VECTOR (7 downto 0);
           hex2  : out STD_LOGIC_VECTOR (7 downto 0);
           hex3  : out STD_LOGIC_VECTOR (7 downto 0));
end lab13_G09;

architecture Behavioral of lab13_G09 is
    signal minute_count : integer range 0 to 59 := 59;
    signal second_count : integer range 0 to 59 := 57;
    signal clk_counter  : integer range 0 to 50000000 := 0; -- Assuming a 50 MHz clock
   
    -- Define the seven-segment codes for numbers 0 through 9
    type segment_array is array (0 to 9) of std_logic_vector(7 downto 0);
    signal segment_codes : segment_array := (
		"01000000",  -- 0
		"01111001",  -- 1
		"00100100",  -- 2
		"00110000",  -- 3
		"00011001",  -- 4
		"00010010",  -- 5
		"00000010",  -- 6
		"01111000",  -- 7
		"00000000",  -- 8
		"00010000"   -- 9
    );

begin
    process(clk)
    begin
        if rising_edge(clk) then
            -- Increment the second count every clock cycle
            if clk_counter = 50000000 then
                clk_counter <= 0;
                if second_count = 59 then
                    second_count <= 0;
                    minute_count <= minute_count + 1;
                    if minute_count = 59 then
                        minute_count <= 0;
                    else
                        minute_count <= minute_count + 1;
                    end if;
                else
                    second_count <= second_count + 1;
                end if;
            else
                clk_counter <= clk_counter + 1;
            end if;
        end if;
    end process;

    -- Output the seven-segment code for the tens and units place of the minutes
    hex3 <= segment_codes(minute_count / 10);
    hex2 <= segment_codes(minute_count mod 10);
   
    -- Output the seven-segment code for the tens and units place of the seconds
    hex1 <= segment_codes(second_count / 10);
    hex0 <= segment_codes(second_count mod 10);

end Behavioral;